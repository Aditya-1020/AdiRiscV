import riscv_pkg::*;

module branch_predictor (
    input logic curr_fetch_pc,
    output branch_pred_t prediction_out;
);

    branch_pred_state_e state, next_state;

    

endmodule