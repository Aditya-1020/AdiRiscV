import riscv_pkg::*;

module wb_stage (

);

    timeunit 1ns;
    timeprecision 1ps;


    


endmodule